module andgate(a, b, Q);
input a, b;
output Q;

assign Q = a & b;

endmodule

